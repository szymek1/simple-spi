`ifndef PARAMS_V
`define PARAMS_V

// PWM (LED control)
`define LED_MIN_BRIGHTNESS 5  // minimal level of brightness in %
`define LED_MAX_BRIGHTNESS 90 // maximal level of brightness in %


`endif // PARAMS_V
