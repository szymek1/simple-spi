//////////////////////////////////////////////////////////////////////////////////
// Company: ISAE
// Engineer: Szymon Bogus
//
// Create Date: 24/07/2025
// Design Name:
// Module Name: spi_master_mock
// Project Name: simple-spi
// Target Devices: Zybo Z7-20
// Tool Versions:
// Description: Mock-up ESP32 SPI Master designed to simulate the micrcontroller
//              SPI master behavior used to validate actually synthesizeable
//              FPGA SPI slave.
//
// Dependencies: params.vh
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns/1ps
`include "../include/params.vh"


module spi_master_mock (

);



endmodule