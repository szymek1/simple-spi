//////////////////////////////////////////////////////////////////////////////////
// Company: ISAE
// Engineer: Szymon Bogus
//
// Create Date: 21/07/2025
// Design Name:
// Module Name: pmw
// Project Name: simple-spi
// Target Devices: Zybo Z7-20
// Tool Versions:
// Description: Pulse-Width-Modulation module. It receives the information what
//              should be the level of a selected LED brightness and outputs
//              control PWM signal.
//
// Dependencies: params.vh
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
`include "../include/params.vh"


module pmw (
    

);
endmodule
