`ifndef PARAMS_V
`define PARAMS_V

// PWM (LED control)
`define BRIGHTNESS_WIDTH   7  // brightness level can vary: 0%-100%; 7-bit number required to store the input value
`define LED_MIN_BRIGHTNESS 5  // minimal level of brightness in %- min. duty cycle
`define LED_MAX_BRIGHTNESS 90 // maximal level of brightness in %- max. duty cycle
`define 


`endif // PARAMS_V
